`define CONNECTAL_MEMORY
`define OUT_OF_ORDER
